library verilog;
use verilog.vl_types.all;
entity CA6_vlg_vec_tst is
end CA6_vlg_vec_tst;
