library verilog;
use verilog.vl_types.all;
entity ca5_vlg_vec_tst is
end ca5_vlg_vec_tst;
